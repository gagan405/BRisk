library IEEE;
library gaisler;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_misc.all;
use IEEE.numeric_std.all;
use work.types.all;
use gaisler.leon3.all;

entity cpu is
	generic (
		CACHE_LINE_ADR  :     natural := 4;
		CACHE_BLOCK_ADR :     natural := 4;
		WRITE_FIFO_ADR  :     natural := 4);
	port (
		clk             : in  std_logic;
		res             : in  std_logic;
		mem_in          : out memory_in;
		mem_out         : in  memory_out;
		irqi            : in  l3_irq_in_type;
		irqo            : out l3_irq_out_type);
end cpu;

architecture structure of cpu is
--signals for IF unit.
signal instr_fetch_mem_out, tie_down : memory_in;-- output memory port of instruction fetch unit connected to input port arbiter.
signal instr_fetch_mem_in  : memory_out; -- output port of arbiter connected to input port of instruction fetch
--signals for memory arbiter
signal wb_memory_in_tb,memory_port_input : memory_in;
signal wb_memory_out_tb,memory_port_output : memory_out;
--signals for testbench
signal ctrl_stall_tb, stall_req_if_tb, branch_tb : std_logic; 
signal branch_target_tb, counter :std_logic_vector(31 downto 0);
signal ins_tb:instruction;
signal decode_out_tb : instruction_decoded;
signal operand_output_tb: operand_type; 
signal memory_out_ldsr_tb: memory_out;
signal write_back_out_tb : write_back;
signal stall_glb_tb,stall_out_if_tb, stall_req_ldsr_tb : std_logic;
signal write_back_input_tb : write_back;
signal decode_out_exe_tb : instruction_decoded; -- decode out from exe unit
signal branch_out_tb : branch; -- beanch out from exe unit
signal store_data_out_tb : std_logic_vector(31 downto 0);
signal exe_out_tb : std_logic_vector(31 downto 0);
signal write_back_ex_tmp : write_back;
signal stall_to_if, stall_to_id, stall_to_ex, stall_to_wb, branch_detect : std_logic;

--signals for cache unit
signal cache_mem_out :  memory_in;
signal cache_mem_in : memory_out;

component mem_arbiter
	port (
        clk: in std_logic;
        res: in std_logic;
        port1_in: in memory_in;
        port2_in: in memory_in;
        port1_out: out memory_out;
        port2_out: out memory_out;
        mem_in: out memory_in;
        mem_out: in memory_out
	);
end component;

component instr_fetch
	port (
	clk: in std_logic;
	ctrl: in control; -- reset and stall control signal input
	stall_req: out std_logic; -- ouput stall control signal generated by instruction fectch unit
	brn : in branch;-- branch control signal and branch address input.
	req_mem: out memory_in; -- memory port connecting to input port of Memory
	rd_mem: in memory_out;  -- port connecting to output port of memory.
	ins: out instruction
	);
end component;

component opcode_disassembler -- used for debugging 
    PORT (Opcode : in Std_Logic_Vector(31 downto 0));
END component;

component instr_decode
	port (
	clk: in std_logic;
	ctrl: in control; 
	ins: in instruction; 
	instrn_decode_out: out instruction_decoded; 
	operand_output: out operand_type;
	branch : 	in  std_logic;
        write_back_ex: in write_back;
	write_back_input: in write_back      
	);
end component;

component instr_exe
	port (
	clk: in std_logic;
	ctrl: in control; --reset and stall inputs
	instruction_decode_in: in instruction_decoded; 
	instruction_decode_out: out instruction_decoded; 
	operand_in: in operand_type; --operand outputs of instrn decode block. 
	branch_out: out branch; --branch control signal and target address.
	exe_out : out std_logic_vector(31 downto 0); --output of the adder.
	wb_in : in write_back;
	write_back_ex: out write_back;
	store_data_out: out Tdata --data to be written to memory is provided in this register.
	);
end component;

component load_store_unit
	port (
	-- control inputs
	clk         :       in std_logic;
	ctrl        :       in control;
	-- outputs 
	stall_req   :       out std_logic;
	wb          :       out write_back;
	-- memory access ports
	to_memory   :       out memory_in;
	from_memory :       in  memory_out;
	-- from the Execution unit
	ins_decoded :       in instruction_decoded;
	data        :       in Tdata;
	addr        :       in Tadr
	);
end component;

component instruction_cache
  generic (
  LINE_ADR : natural := 4; --no of bits for line address
  BLOCK_ADR : natural := 4 -- no of bits for block address for each line.
  );
  
  port (
    clk : in std_logic;
    res : in std_logic;
    
    cpu_from : in memory_in;
    cpu_to   : out memory_out;
    memory_to   : out memory_in;
    memory_from : in memory_out
  );
end component;

begin
	tie_down.enable <= '0';
	tie_down.adr <= (others => '0');
	tie_down.data <= (others => '0');
	tie_down.we <= '0';

	mem_in <= memory_port_input;
	memory_port_output <= mem_out;
	
	write_back_input_tb.d <= (others => '0');
	write_back_input_tb.idx_d <= (others => '0');
	write_back_input_tb.d_valid <= '0';
	ctrl_stall_tb <= '0';

	stall_to_if <= stall_req_ldsr_tb;
        stall_to_id <= stall_out_if_tb or stall_req_ldsr_tb;--stall_out_if_tb; --
	stall_to_ex <= stall_out_if_tb or stall_req_ldsr_tb;--stall_out_if_tb; --
	stall_to_wb <= stall_out_if_tb;
	branch_detect <= branch_out_tb.branch;


	mem_arb:mem_arbiter
	port map (
		clk => clk,
		res => res,
		port1_in =>cache_mem_out,  --instr_fetch_mem_out,
		port2_in => wb_memory_in_tb,	
		port1_out =>cache_mem_in,  --instr_fetch_mem_in ,
		port2_out => wb_memory_out_tb,	--
		mem_in => memory_port_input,
		mem_out=> memory_port_output
		);

        instruction_fetch:instr_fetch
	port map (
		clk => clk,
		ctrl.res => res,
		ctrl.stall => stall_to_if,
		stall_req => stall_out_if_tb, 
--		brn.branch => branch_tb,
--		brn.target => branch_target_tb,
		brn => branch_out_tb,
		req_mem=>instr_fetch_mem_out,
		rd_mem => instr_fetch_mem_in,
		ins => ins_tb
		);

	opcode_dis:opcode_disassembler
	port map (
		Opcode => ins_tb.ir
		);

	instruction_decode:instr_decode
	port map (
		clk => clk,
		ctrl.res => res,
		ctrl.stall => stall_to_id,
		ins => ins_tb,
		branch => branch_detect,
		instrn_decode_out => decode_out_tb,
		operand_output => operand_output_tb,
		write_back_ex => write_back_ex_tmp,
		write_back_input => write_back_out_tb
		);

	instruction_execute:instr_exe
	port map (
		clk => clk,
		ctrl.res => res,
		ctrl.stall => stall_to_ex,
		instruction_decode_in => decode_out_tb,
		instruction_decode_out => decode_out_exe_tb,
		operand_in => operand_output_tb,
		branch_out => branch_out_tb,
		wb_in => write_back_out_tb,
		write_back_ex => write_back_ex_tmp,
		exe_out => exe_out_tb,
		store_data_out =>store_data_out_tb
		);

	instruction_load_store:load_store_unit
	port map(
		-- control inputs
		clk => clk,
		ctrl.res => res,
		ctrl.stall => stall_to_wb,
		-- outputs 
		stall_req  => stall_req_ldsr_tb,
		wb  => write_back_out_tb,
		-- memory access ports
		to_memory  => wb_memory_in_tb,
		from_memory  => wb_memory_out_tb,
		-- from the Execution unit
		ins_decoded  => decode_out_exe_tb,
		data  =>store_data_out_tb,
		addr => exe_out_tb
		);

	instruction_cache_unit: instruction_cache
	generic map (
		LINE_ADR =>  CACHE_LINE_ADR, --no of bits for line address
		BLOCK_ADR => CACHE_BLOCK_ADR -- no of bits for block address for each line.
		)
	port map (
		clk  => clk,
		res  => res,
		cpu_from => instr_fetch_mem_out,
		cpu_to => instr_fetch_mem_in,
		memory_to   => cache_mem_out,
		memory_from => cache_mem_in
		);


--	stall_check: process (clk)
--	begin
--	  if (clk'event and clk = '1') then
--		  if (res = '1') then
--			ctrl_stall_tb <= '0';
--			counter <= (others => '0');
--		  else
--			counter <= std_logic_vector(unsigned(counter)+1);
--			if (counter = x"00000002") then
--			   ctrl_stall_tb <= '1';
--			elsif (counter = x"00000003") then
--			   ctrl_stall_tb <= '1';
--			elsif (counter = x"00000004") then
--			   ctrl_stall_tb <= '1';
--			elsif (counter = x"00000005") then
--			   ctrl_stall_tb <= '1';
--			elsif (counter = x"00000008") then
--			   ctrl_stall_tb <= '1';
--			elsif (counter = x"00000009") then
--			   ctrl_stall_tb <= '0';
--			elsif (counter = x"0000000a") then
--			   ctrl_stall_tb <= '1';
--			  else 
--			   ctrl_stall_tb <= '0';
--			end if;
--		  end if;
--	  end if;
--	end process;
--
	branch_check: process (clk)
	begin
	  if (clk'event and clk = '1') then
		  if (res = '1') then
			branch_tb <= '0';
			branch_target_tb <= (others => '0');
		  end if;
	   end if;
	end process;

end structure;
